<glayout.spice.netlist.Netlist object at 0x72ecfd7a30a0>