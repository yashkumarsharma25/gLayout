<glayout.spice.netlist.Netlist object at 0x752bbbe37910>